/*
 * Module: MVAU Streaming Block (mvau_stream.sv)
 * 
 * Author(s): Syed Asad Alam <syed.asad.alam@tcd.ie>
 * 
 * This file lists an RTL implementation of the matrix-vector multiplication unit
 * based on streaming weights. It can either be part of the Matrix-Vector-Activation Unit
 * or run independently
 *
 * This material is based upon work supported, in part, by Science Foundation
 * Ireland, www.sfi.ie under Grant No. 13/RC/2094 and, in part, by the 
 * European Union's Horizon 2020 research and innovation programme under the 
 * Marie Sklodowska-Curie grant agreement Grant No.754489. 
 * 
 * Inputs:
 * aresetn - Active low, synchronous reset
 * aclk - Main clock
 * rready - Input ready
 * in_v - Input valid when input activation is valid
 * [TI-1:0] in_act - Input activation stream, word length TI=TSrcI*SIMD
 * in_wgt_v - Input weight valid
 * [0:SIMD*TW-1:0] in_wgt [0:PE-1] - Input weight stream
 * 
 * Outputs:			       
 * wready - Output ready
 * wmem_ready - Output ready for weight 
 * out_v        - Output stream valid
 * [TO-1:0] out - Output stream, word length TO=TDstI*PE
 * 
 * Parameters:
 * KDim         - Kernel dimensions                                                                    
 * IFMCh        - Input feature map channels                                                           
 * OFMCh        - Output feature map channels or the number of filter banks                            
 * IFMDim       - Input feature map dimensions                                                       
 * PAD          - Padding around the input feature map                                                  
 * STRIDE       - Number of pixels to move across when applying the filter                           
 * OFMDim       - Output feature map dimensions                                                      
 * MatrixW      - Width of the input matrix                                                         
 * MatrixH      - Heigth of the input matrix                                                        
 * SIMD         - Number of input columns computed in parallel                                         
 * PE           - Number of output rows computed in parallel                                             
 * WMEM_DEPTH   - Depth of each weight memory                                                    
 * MMV          - Number of output pixels computed in parallel                                          
 * TSrcI        - DataType of the input activation (as used in the MAC)                               
 * TSrcI_BIN    - Indicates whether the 1-bit TSrcI is to be interpreted as special +1/-1 or not
 * TI           - SIMD times the word length of input stream                                             
 * TW           - Word length of individual weights                                                      
 * TW_BIN       - Indicates whether the 1-bit TW is to be interpreted as special +1/-1 or not      
 * TDstI        - DataType of the output activation (as generated by the activation)                  
 * TO           - PE times the word length of output stream                                             
 * TA           - PE times the word length of the activation class (e.g thresholds)                     
 * USE_DSP      - Use DSP blocks or LUTs for MAC                                                    
 * MVAU_STREAM  - Top module is not MVAU Stream                                                 
 * USE_ACT      - Use activation after matrix-vector activation       
 * SF=MatrixW/SIMD - Number of vertical weight matrix chunks and depth of the input buffer
 * NF=MatrixH/PE   - Number of horizontal weight matrix chunks
 * SF_T            - log_2(SF), determines the number of address bits for the input buffer
 * NF_T            - log_2(NF), word length of the NF counter to control reading and writing from the input buffer
 * */

`timescale 1ns/1ns

module mvau_stream #(
		     parameter int KDim=2, // Kernel dimensions
		     parameter int IFMCh=2,// Input feature map channels
		     parameter int OFMCh=2,// Output feature map channels or the number of filter banks
		     parameter int IFMDim=2, // Input feature map dimensions
		     parameter int PAD=0, // Padding around the input feature map
		     parameter int STRIDE=1, // Number of pixels to move across when applying the filter
		     parameter int OFMDim=1, // Output feature map dimensions
		     parameter int MatrixW=8, // Width of the input matrix
		     parameter int MatrixH=2, // Heigth of the input matrix
		     parameter int SIMD=2, // Number of input columns computed in parallel
		     parameter int PE=2, // Number of output rows computed in parallel
		     parameter int WMEM_DEPTH=4, // Depth of each weight memory
		     parameter int MMV=1, // Number of output pixels computed in parallel
		     parameter int TSrcI=4, // DataType of the input activation (as used in the MAC)
		     parameter int TSrcI_BIN = 0, // Indicates whether the 1-bit TSrcI is to be interpreted as special +1/-1 or not
		     parameter int TI=8, // SIMD times the word length of input stream
		     parameter int TW=1, // Word length of individual weights
		     parameter int TW_BIN = 0, // Indicates whether the 1-bit TW is to be interpreted as special +1/-1 or not
		     parameter int TDstI=8, // DataType of the output activation (as generated by the activation) 
		     parameter int TO=16, // PE times the word length of output stream   
		     parameter int TA=16, // PE times the word length of the activation class (e.g thresholds)
		     parameter int USE_DSP=0, // Use DSP blocks or LUTs for MAC
		     parameter int MVAU_STREAM=1, // Top module is not MVAU Stream
		     parameter int USE_ACT=0)     // Use activation after matrix-vector activation	      
   (
    input logic 		 aresetn,
    input logic 		 aclk,
    input logic 		 rready,
    output logic 		 wready,
    output logic 		 wmem_wready,
    input logic 		 in_v,
    input logic [TI-1:0] 	 in_act ,
    input logic 		 in_wgt_v, // Input valid from the weight stream
    input logic [0:PE*SIMD*TW-1] in_wgt, // Streaming weight tile
    output logic 		 out_v, // Ouptut valid
    output logic [TO-1:0] 	 out);

   /*
    * Local parameters
    * */
   // Parameter: SF
   // Number of vertical matrix chunks to be processed in parallel by one PE
   localparam int SF=MatrixW/SIMD; // Number of vertical matrix chunks
   // Parameter: NF
   // Number of horizontal matrix chunks to be processed by PEs in parallel
   localparam int NF=MatrixH/PE; // Number of horizontal matrix chunks
   // Parameter: SF_T
   // Address word length of the buffer
   localparam int SF_T=$clog2(SF); // Address word length for the input buffer
   // Parameter: NF_T
   // Word length of the NF counter to control reading and writing from the input buffer
   localparam int 	    NF_T=$clog2(NF); // For nf_cnt	 
   
   /**
    * Internal Signals
    * **/
   // Signal: in_act_reg
   // Input activation stream synchronized to clock
   logic [TI-1:0] 		       in_act_reg;
   // Signal: in_wgt_reg
   // Streaming weight tile synchronized to clock
   logic [0:SIMD-1][TW-1:0] 	       in_wgt_reg [0:PE-1];
   // Internal signals for the input buffer and the control block
   // Signal: ib_wen
   // Write enable for the input buffer
   logic 		      ib_wen;
   // Signal: ib_ren
   // Read enable for the input buffer
   logic 		      ib_ren;
   // Signal: sf_clr
   // Resets the accumulator as well the sf_cnt
   logic 		      sf_clr;
   // Signal out_act
   // Output of the input buffer
   logic [TI-1:0] 	      out_act;    
   // Signal: out_pe
   // Holds the output from parallel PEs
   logic [0:PE-1][TDstI-1:0]  out_pe;
   // Signal: out_pe_v
   // Output valid signal from each PE
   logic [0:PE-1] 	      out_pe_v;
   // Signal: do_mvau_stream   
   // Controls how long the MVAU operation continues
   // Case 1: NF=1 => do_mvau_stream = in_v (input buffer not reused)
   // Case 2: NF>1 => do_mvau_stream = in_v | (~(nf_clr&sf_clr)) (input buffer reused)
   logic 		      do_mvau_stream;
   // Signal: in_wgt2d
   // Copy of input weight stream with packed and  unpacked dimension
   logic [0:SIMD*TW-1] 	      in_wgt2d [0:PE-1];
   // Signal: wait_rready
   // Indicates that the design is waiting for ready after valid is asserted
   logic 		      wait_rready;
   

   // Always_FF: DO_MVAU_STREAM
   // Registered signal indicating when to perform the
   // Matrix vector multiplication
   // Dependent on valids and readys
   always_ff @(posedge aclk) begin
      if(!aresetn) 
	do_mvau_stream <= 1'b0;
      else
	do_mvau_stream <= in_v & wready | in_wgt_v & wmem_wready;
   end
   
   // Copying the packed input weight array
   // to packed/unpacked array
   generate
      for(genvar p = 0; p < PE; p++) begin
	 assign in_wgt2d[p] = in_wgt[SIMD*TW*p:SIMD*TW*p+(SIMD*TW-1)];	 
      end
   endgenerate

   // Only registering weights
   // when the stream unit is the top level unit
   generate
      if(MVAU_STREAM==1) begin: MVAU_STREAM_TOP
   	 // Always_FF: WGT_REG
   	 // Register the input weight stream
	 // Only when the stream unit is the top level unit
   	 always_ff @(posedge aclk) begin
   	    if(!aresetn) begin
   	       for(int i = 0; i < PE; i++)
   		 in_wgt_reg[i] <= 'd0;
   	    end
   	    else begin
   	       for(int i = 0; i < PE; i++)
   		 in_wgt_reg[i] <= in_wgt2d[i];
   	    end
   	 end
      end // block: MVAU_STREAM_TOP      
      else begin: MVAU_BATCH_TOP
	 always_comb begin
	    for(int i = 0; i < PE; i++)
	      in_wgt_reg[i] = in_wgt2d[i];
	 end	 
      end      
   endgenerate
   assign in_act_reg = in_act;

   // Always_FF: WAIT_READY
   // Indicates if after assertion of output valid,
   // input ready is not asserted to read the output
   // Helps in pausing all computations until the output is consumed
   always_ff @(posedge aclk) begin
      if(!aresetn)
	wait_rready <= 1'b0;
      else if(rready)
	wait_rready <= 1'b0;
      else if(out_v)
	wait_rready <= 1'b1;
   end
      
   /*
    * Control logic for reading and writing to input buffer
    * and the input buffer itself
    * Four cases:
    * Case 1: SF=1, NF=1
    * Case 2: SF=1, NF>1
    * Case 3: SF>1, NF=1
    * Case 4: SF=1, NF=1
    * */
   if(SF==1) begin: SF_1
      if(NF==1) begin: NF_1
	 // Signal: sf_cnt
	 // Counter keeping track of SF and also address to input buffer
	 // One bit in case SF=1
	 // log2(SF) bits otherwise
	 logic sf_cnt;
	 mvau_stream_control_block #(
				     .SF(SF),
				     .NF(NF),
				     .SF_T(1),
				     .NF_T(1)
				     )
	 mvau_stream_cb_inst (.aresetn,
			      .aclk,
			      .in_v(in_v),
			      .ib_wen,
			      .ib_ren,
			      .wait_rready,
			      .wready,
			      .wmem_wready,
			      .sf_clr,
			      .sf_cnt);
	 mvau_inp_buffer #(
			   .TI(TI),
			   .BUF_LEN(SF),
			   .BUF_ADDR(1))
	 mvau_inb_inst (
			.aclk,
			.aresetn,
			.in(in_act_reg),
			.wr_en(ib_wen),
			.rd_en(ib_ren),
			.addr(sf_cnt),
			.out(out_act));
      end // block: NF_1      
      else begin: NF_N
	 logic sf_cnt;
	 mvau_stream_control_block #(
				     .SF(SF),
				     .NF(NF),
				     .SF_T(1),
				     .NF_T(NF_T)
				     )
	 mvau_stream_cb_inst (.aresetn,
			      .aclk,
			      .in_v(in_v),
			      .ib_wen,
			      .ib_ren,
			      .wait_rready,
			      .wready,
			      .wmem_wready,
			      .sf_clr,
			      .sf_cnt);
	 mvau_inp_buffer #(
			   .TI(TI),
			   .BUF_LEN(SF),
			   .BUF_ADDR(1))
	 mvau_inb_inst (
			.aclk,
			.aresetn,
			.in(in_act_reg),
			.wr_en(ib_wen),
			.rd_en(ib_ren),
			.addr(sf_cnt),
			.out(out_act));
      end // block: NF_N
   end // block: SF_1   
   else begin: SF_N
      if(NF==1) begin: NF_1	 
	 logic [SF_T-1:0] 	      sf_cnt;
	 mvau_stream_control_block #(
				     .SF(SF),
				     .NF(NF),
				     .SF_T(SF_T),
				     .NF_T(1)
				     )
	 mvau_stream_cb_inst (.aresetn,
			      .aclk,
			      .in_v(in_v),
			      .ib_wen,
			      .ib_ren,
			      .wait_rready,
			      .wready,
			      .wmem_wready,
			      .sf_clr,
			      .sf_cnt);
	  mvau_inp_buffer #(
			   .TI(TI),
			   .BUF_LEN(SF),
			   .BUF_ADDR(SF_T))
	 mvau_inb_inst (
			.aclk,
			.aresetn,
			.in(in_act_reg),
			.wr_en(ib_wen),
			.rd_en(ib_ren),
			.addr(sf_cnt),
			.out(out_act));
      end // block: NF_1
      else begin: NF_N
	 logic [SF_T-1:0] 	      sf_cnt;
	 mvau_stream_control_block #(
				     .SF(SF),
				     .NF(NF),
				     .SF_T(SF_T),
				     .NF_T(NF_T)
				     )
	 mvau_stream_cb_inst (.aresetn,
			      .aclk,
			      .in_v(in_v),
			      .ib_wen,
			      .ib_ren,
			      .wait_rready,
			      .wready,
			      .wmem_wready,
			      .sf_clr,
			      .sf_cnt);
	  mvau_inp_buffer #(
			   .TI(TI),
			   .BUF_LEN(SF),
			   .BUF_ADDR(SF_T))
	 mvau_inb_inst (
			.aclk,
			.aresetn,
			.in(in_act_reg),
			.wr_en(ib_wen),
			.rd_en(ib_ren),
			.addr(sf_cnt),
			.out(out_act));
      end // block: NF_N
   end // block: SF_N
      
   
   /**
    * Generating instantiations of all processing elements
    * Each PE reads in different set of weights
    * Each PE reads in the same set of activation
    * Each PE outputs TDstI bits
    * Output of each PE packed into one array of size TO
    * */
   generate
      for(genvar pe_ind = 0; pe_ind < PE; pe_ind = pe_ind+1)
	begin: PE_GEN
	   mvu_pe #(
		    .SIMD(SIMD),
		    .PE(PE),
		    .TSrcI(TSrcI),
		    .TSrcI_BIN(TSrcI_BIN),
		    .TI(TI),
		    .TW(TW),
		    .TW_BIN(TW_BIN),
		    .TDstI(TDstI),
		    .TO(TO))
	   mvu_pe_inst( // Mapping the I/O blocks
			.aresetn,
			.aclk,
			.sf_clr,
			.do_mvau_stream,
			.in_act(out_act),
			.in_wgt(in_wgt_reg[pe_ind]),
			.out_v(out_pe_v[PE-pe_ind-1]),
			.out(out_pe[PE-pe_ind-1]) // Each PE contribution TDstI bits in the output
			);
	end
   endgenerate

   // A place holder for the activation unit to be implemented later
   if(USE_ACT==1) begin: ACT
   end
   else begin: NO_ACT
      // Two cases handled here
      // Case 1: MVAU Stream unit is top level DUT
      // Case 2: MVAU Stream unit is not top level DUT
      if(MVAU_STREAM==1) begin: MVAU_STREAM_OUT
	 // Case 1: MVAU Stream unit is top level DUT
	 logic out_pe_v_one;
	 assign out_pe_v_one = |out_pe_v;

	 logic out_pe_valid_hold;
	 logic [TO-1:0] out_pe_hold;
	 
	 // Always_FF: OUT_STREAM_V_HOLD
	 // Saving the 2nd PE valid if it comes
	 // before previous output consumed by the slave interface
	 always_ff @(posedge aclk) begin
	    if(!aresetn)
	      out_pe_valid_hold <= 1'b0;
	    else if(~out_v & out_pe_valid_hold) // Finish hold
	      out_pe_valid_hold <= 1'b0;
	    else if(out_pe_v_one & out_v) // Start hold
	      out_pe_valid_hold <= 1'b1;	    
	 end

	 // Always_FF: OUT_PE_HOLD
	 // Saving the 2nd PE output if it comes
	 // before previous output consumed by the slave interface
	 always_ff @(posedge aclk) begin
	    if(!aresetn)
	      out_pe_hold <= 'd0;
	    else if(out_pe_v_one & out_v) // Start hold
	      out_pe_hold <= out_pe;
	 end	 

	 // Always_FF: OUT_PE_REG
	 // Registering the output activation stream
	 // Three cases
	 // a) Hold output if input ready not asserted
	 // b) Read PE output
	 // c) Read the saved PE output
	 always_ff @(posedge aclk) begin
	    if(!aresetn)
	      out <= 'd0;
	    else if(out_v & ~rready)
	      out <= out;
	    else if(out_pe_v_one)
	      out <= out_pe;
	    else if(out_pe_valid_hold)
	      out <= out_pe_hold;	    
	 end
	 // Always_FF: OUT_V_REG
	 // Registering the output activation stream valid signal
	 // Asserted when either there is an ouptut asserted by the PEs
	 // or an output held due to non-consumption
	 // When output is consumed, as shown by an asserted ready input signal,
	 // output valid is deasserted
	 always_ff @(posedge aclk) begin
	    if(!aresetn) 
	      out_v <= 1'b0;	    	    
	    else if(out_pe_v_one)
	      out_v <= 1'b1;
	    else if(out_v & rready)
	      out_v <= 1'b0;	    
	    else if(out_pe_valid_hold)
	      out_v <= 1'b1;	    
	 end
      end // block: MVAU_STREAM_OUT
      else begin: MVAU_BATCH_OUT
	 // Case 2: MVAU Stream is not top level DUT
	 // Simply passing the outputs to the Batch unit
	 assign out_v = (|out_pe_v);
	 assign out = out_pe;
      end
   end // block: NO_ACT
   
endmodule // mvau_stream
