/*********************************************/
/*********************************************/
/*** Package for definitions and constants ***/
/*** for multiply-vector activation unit   ***/
/*********************************************/
/*********************************************/

/**
 * Defines the following parameters
 * that control the generation of 
 * the matrix vector activation unit
 * 
 * VERION
 * KDim                                // Kernel dimensions                                                             
 * IFMCh                               // Input feature map channels                                                    
 * OFMCh                               // Output feature map channels                                                   
 * IFMDim		               // Input feature map dimensions                                                
 * PAD                                 // Padding around the input feature map                     
 * STRIDE		               // Number of pixels to move across when applying the filter 
 * OFMDim=(IFMDim-KDim+2*PAD)/STRIDE+1 // Output feature map dimensions                                               
 * MatrixW=KDim*KDim*IFMCh             // Width of the input matrix                                  
 * MatrixH=OFMCh                       // Heigth of the input matrix                                             
 * SIMD                                // Number of input columns computed in parallel                                 
 * PE                                  // Number of output rows computed in parallel                                      
 * MMV                                 // Number of output pixels computed in parallel                                   
 * TSrcI                               // DataType of the input activation (as used in the MAC)                        
 * TDstI                               // DataType of the output activation (as generated by the activation)           
 * TWeightI                            // DataType of the weights and how to access them in the array (Class in HLS)
 * TI                                  // SIMD times the word length of input stream                                      
 * TO                                  // PE times the word length of output stream                                      
 * TW                                  // Word length of individual weights                                               
 * TA                                  // PE times the word length of the activation class (e.g thresholds)              
 * USE_DSP                             // Use DSP blocks or LUTs for MAC (future extension)                                       
 * INST_WMEM                           // Instantiate weight memory; if needed
 * USE_ACT                             // Use activation after matrix-vector activation
 * **/

`ifndef MVAU_DEFN_PKG // if the already-compiled flag is not set
 `define MVAU_DEFN_PKG //set the flag
package mvau_defn;
   parameter VERSION = "0.1";
   parameter int KDim=5; // Kernel dimensions
   parameter int IFMCh=3;// Input feature map channels
   parameter int OFMCh=8;// Output feature map channels or the number of filter banks
   parameter int IFMDim=32; // Input feature map dimensions
   parameter int PAD=0;    // Padding around the input feature map
   parameter int STRIDE=1; // Number of pixels to move across when applying the filter
   parameter int OFMDim=(IFMDim-KDim+2*PAD)/STRIDE+1; // Output feature map dimensions
   parameter int MatrixW=KDim*KDim*IFMCh;   // Width of the input matrix                                          
   parameter int MatrixH=OFMCh; // Heigth of the input matrix   
   parameter int SIMD=5; // Number of input columns computed in parallel                       
   parameter int PE=4; // Number of output rows computed in parallel                         
   parameter int WMEM_DEPTH=(KDim*KDim*IFMCh*OFMCh)/(SIMD*PE); // Depth of each weight memory   
   parameter int MMV=1; // Number of output pixels computed in parallel                       
   parameter int TSrcI=4; // DataType of the input activation (as used in the MAC)   
   parameter int TI=SIMD*TSrcI; // SIMD times the word length of input stream
   parameter int TWeightI=1; // DataType of the weights and how to access them in the array (Class in HLS)
   parameter int TW=4; // Word length of individual weights   
   parameter int TDstI=4; // DataType of the output activation (as generated by the activation) 
   parameter int TO=PE*TDstI; // PE times the word length of output stream   
   parameter int TA=16; // PE times the word length of the activation class (e.g thresholds)
   parameter int USE_DSP=0; // Use DSP blocks or LUTs for MAC
   parameter int INST_WMEM=0; // Instantiate weight memory; if needed
   parameter int USE_ACT=0;     // Use activation after matrix-vector activation
   
endpackage
   
   import mvau_defn::*; // import package into $unit compilation space
`endif

