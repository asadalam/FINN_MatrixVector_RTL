/*********************************************/
/*********************************************/
/*** Package for definitions and constants ***/
/*** for multiply-vector activation unit   ***/
/*********************************************/
/*********************************************/

`ifndef MVAU_DEFN_PKG // if the already-compiled flag is not set
 `define MVAU_DEFN_PKG //set the flag
package mvau_defn;
   parameter VERSION = "0.1";
   parameter int KDim=2; // Kernel dimensions
   parameter int IFMCh=4;// Input feature map channels
   parameter int OFMCh=4;// Output feature map channels
   parameter int IFMDim=4; // Input feature map dimensions
   parameter int OFMDim=3; // Output feature map dimensions
   parameter int MatrixW=KDim*KDim*IFMCh;   // Width of the input matrix                                          
   parameter int MatrixH=OFMCh; // Heigth of the input matrix
   parameter int SIMD=2; // Number of input columns computed in parallel                       
   parameter int PE=2; // Number of output rows computed in parallel                         
   parameter int MMV=1; // Number of output pixels computed in parallel                       
   parameter int TSrcI=1; // DataType of the input activation (as used in the MAC)              
   parameter int TDstI=1; // DataType of the output activation (as generated by the activation) 
   parameter int TWeightI=1; // DataType of the weights and how to access them in the array
   parameter int TI=2; // SIMD times the word length of input stream
   parameter int TO=2; // PE times the word length of output stream
   parameter int TW=2; // SIMD times the word length of weight stream
   parameter int TA=2; // PE times the word length of the activation class (e.g thresholds)
   parameter int USE_DSP=0; // Use DSP blocks or LUTs for MAC
   parameter int INST_WMEM=0; // Instantiate weight memory; if needed
   parameter int USE_ACT=0;     // Use activation after matrix-vector activation
   localparam int SF=MatrixW/SIMD; // Number of vertical matrix chunks
   localparam int NF=MatrixH/PE; // Number of horizontal matrix chunks
   localparam int SF_T=$clog2(SF); // Address word length for the input buffer
endpackage
   
   import mvau_defn::*; // import package into $unit compilation space
`endif

